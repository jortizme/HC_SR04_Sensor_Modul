# Input signal von außen mussen hier synchrnoiwist werden